VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_1024x32_upper
  FOREIGN fakeram45_1024x32_upper 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 152.190 BY 107.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 12.880 0.070 12.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 14.560 0.070 14.630 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 16.240 0.070 16.310 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 17.920 0.070 17.990 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 21.280 0.070 21.350 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 37.240 0.070 37.310 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 38.080 0.070 38.150 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 38.920 0.070 38.990 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 39.760 0.070 39.830 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 40.600 0.070 40.670 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 42.280 0.070 42.350 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 43.120 0.070 43.190 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 43.960 0.070 44.030 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 45.640 0.070 45.710 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 46.480 0.070 46.550 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 47.320 0.070 47.390 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 51.520 0.070 51.590 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 52.360 0.070 52.430 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 54.040 0.070 54.110 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 54.880 0.070 54.950 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 55.720 0.070 55.790 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 56.560 0.070 56.630 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 57.400 0.070 57.470 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 59.920 0.070 59.990 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 60.760 0.070 60.830 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 61.600 0.070 61.670 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 62.440 0.070 62.510 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 63.280 0.070 63.350 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 64.120 0.070 64.190 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 64.960 0.070 65.030 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 65.800 0.070 65.870 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 66.640 0.070 66.710 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 67.480 0.070 67.550 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 68.320 0.070 68.390 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 69.160 0.070 69.230 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 70.000 0.070 70.070 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 70.840 0.070 70.910 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 71.680 0.070 71.750 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 72.520 0.070 72.590 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 73.360 0.070 73.430 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 74.200 0.070 74.270 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 75.040 0.070 75.110 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 75.880 0.070 75.950 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 76.720 0.070 76.790 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 77.560 0.070 77.630 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 78.400 0.070 78.470 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 79.240 0.070 79.310 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 80.080 0.070 80.150 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 80.920 0.070 80.990 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 81.760 0.070 81.830 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 82.600 0.070 82.670 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 83.440 0.070 83.510 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 84.280 0.070 84.350 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 85.120 0.070 85.190 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 85.960 0.070 86.030 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 88.480 0.070 88.550 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 89.320 0.070 89.390 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 90.160 0.070 90.230 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 91.000 0.070 91.070 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 91.840 0.070 91.910 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 92.680 0.070 92.750 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 93.520 0.070 93.590 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 94.360 0.070 94.430 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 95.200 0.070 95.270 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 96.040 0.070 96.110 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 98.560 0.070 98.630 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 99.400 0.070 99.470 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M18 ;
      RECT 0.000 100.240 0.070 100.310 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M17 ;
      RECT 2.660 2.800 2.940 105.000 ;
      RECT 7.140 2.800 7.420 105.000 ;
      RECT 11.620 2.800 11.900 105.000 ;
      RECT 16.100 2.800 16.380 105.000 ;
      RECT 20.580 2.800 20.860 105.000 ;
      RECT 25.060 2.800 25.340 105.000 ;
      RECT 29.540 2.800 29.820 105.000 ;
      RECT 34.020 2.800 34.300 105.000 ;
      RECT 38.500 2.800 38.780 105.000 ;
      RECT 42.980 2.800 43.260 105.000 ;
      RECT 47.460 2.800 47.740 105.000 ;
      RECT 51.940 2.800 52.220 105.000 ;
      RECT 56.420 2.800 56.700 105.000 ;
      RECT 60.900 2.800 61.180 105.000 ;
      RECT 65.380 2.800 65.660 105.000 ;
      RECT 69.860 2.800 70.140 105.000 ;
      RECT 74.340 2.800 74.620 105.000 ;
      RECT 78.820 2.800 79.100 105.000 ;
      RECT 83.300 2.800 83.580 105.000 ;
      RECT 87.780 2.800 88.060 105.000 ;
      RECT 92.260 2.800 92.540 105.000 ;
      RECT 96.740 2.800 97.020 105.000 ;
      RECT 101.220 2.800 101.500 105.000 ;
      RECT 105.700 2.800 105.980 105.000 ;
      RECT 110.180 2.800 110.460 105.000 ;
      RECT 114.660 2.800 114.940 105.000 ;
      RECT 119.140 2.800 119.420 105.000 ;
      RECT 123.620 2.800 123.900 105.000 ;
      RECT 128.100 2.800 128.380 105.000 ;
      RECT 132.580 2.800 132.860 105.000 ;
      RECT 137.060 2.800 137.340 105.000 ;
      RECT 141.540 2.800 141.820 105.000 ;
      RECT 146.020 2.800 146.300 105.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M17 ;
      RECT 4.900 2.800 5.180 105.000 ;
      RECT 9.380 2.800 9.660 105.000 ;
      RECT 13.860 2.800 14.140 105.000 ;
      RECT 18.340 2.800 18.620 105.000 ;
      RECT 22.820 2.800 23.100 105.000 ;
      RECT 27.300 2.800 27.580 105.000 ;
      RECT 31.780 2.800 32.060 105.000 ;
      RECT 36.260 2.800 36.540 105.000 ;
      RECT 40.740 2.800 41.020 105.000 ;
      RECT 45.220 2.800 45.500 105.000 ;
      RECT 49.700 2.800 49.980 105.000 ;
      RECT 54.180 2.800 54.460 105.000 ;
      RECT 58.660 2.800 58.940 105.000 ;
      RECT 63.140 2.800 63.420 105.000 ;
      RECT 67.620 2.800 67.900 105.000 ;
      RECT 72.100 2.800 72.380 105.000 ;
      RECT 76.580 2.800 76.860 105.000 ;
      RECT 81.060 2.800 81.340 105.000 ;
      RECT 85.540 2.800 85.820 105.000 ;
      RECT 90.020 2.800 90.300 105.000 ;
      RECT 94.500 2.800 94.780 105.000 ;
      RECT 98.980 2.800 99.260 105.000 ;
      RECT 103.460 2.800 103.740 105.000 ;
      RECT 107.940 2.800 108.220 105.000 ;
      RECT 112.420 2.800 112.700 105.000 ;
      RECT 116.900 2.800 117.180 105.000 ;
      RECT 121.380 2.800 121.660 105.000 ;
      RECT 125.860 2.800 126.140 105.000 ;
      RECT 130.340 2.800 130.620 105.000 ;
      RECT 134.820 2.800 135.100 105.000 ;
      RECT 139.300 2.800 139.580 105.000 ;
      RECT 143.780 2.800 144.060 105.000 ;
      RECT 148.260 2.800 148.540 105.000 ;
    END
  END VDD
  OBS
    LAYER M1_m ;
    RECT 0 0 152.190 107.800 ;
    LAYER M19 ;
    RECT 0 0 152.190 107.800 ;
    LAYER M18 ;
    RECT 0.070 0 152.190 107.800 ;
    RECT 0 0.000 0.070 2.800 ;
    RECT 0 2.870 0.070 3.640 ;
    RECT 0 3.710 0.070 4.480 ;
    RECT 0 4.550 0.070 5.320 ;
    RECT 0 5.390 0.070 6.160 ;
    RECT 0 6.230 0.070 7.000 ;
    RECT 0 7.070 0.070 7.840 ;
    RECT 0 7.910 0.070 8.680 ;
    RECT 0 8.750 0.070 9.520 ;
    RECT 0 9.590 0.070 10.360 ;
    RECT 0 10.430 0.070 11.200 ;
    RECT 0 11.270 0.070 12.040 ;
    RECT 0 12.110 0.070 12.880 ;
    RECT 0 12.950 0.070 13.720 ;
    RECT 0 13.790 0.070 14.560 ;
    RECT 0 14.630 0.070 15.400 ;
    RECT 0 15.470 0.070 16.240 ;
    RECT 0 16.310 0.070 17.080 ;
    RECT 0 17.150 0.070 17.920 ;
    RECT 0 17.990 0.070 18.760 ;
    RECT 0 18.830 0.070 19.600 ;
    RECT 0 19.670 0.070 20.440 ;
    RECT 0 20.510 0.070 21.280 ;
    RECT 0 21.350 0.070 22.120 ;
    RECT 0 22.190 0.070 22.960 ;
    RECT 0 23.030 0.070 23.800 ;
    RECT 0 23.870 0.070 24.640 ;
    RECT 0 24.710 0.070 25.480 ;
    RECT 0 25.550 0.070 26.320 ;
    RECT 0 26.390 0.070 27.160 ;
    RECT 0 27.230 0.070 28.000 ;
    RECT 0 28.070 0.070 28.840 ;
    RECT 0 28.910 0.070 31.360 ;
    RECT 0 31.430 0.070 32.200 ;
    RECT 0 32.270 0.070 33.040 ;
    RECT 0 33.110 0.070 33.880 ;
    RECT 0 33.950 0.070 34.720 ;
    RECT 0 34.790 0.070 35.560 ;
    RECT 0 35.630 0.070 36.400 ;
    RECT 0 36.470 0.070 37.240 ;
    RECT 0 37.310 0.070 38.080 ;
    RECT 0 38.150 0.070 38.920 ;
    RECT 0 38.990 0.070 39.760 ;
    RECT 0 39.830 0.070 40.600 ;
    RECT 0 40.670 0.070 41.440 ;
    RECT 0 41.510 0.070 42.280 ;
    RECT 0 42.350 0.070 43.120 ;
    RECT 0 43.190 0.070 43.960 ;
    RECT 0 44.030 0.070 44.800 ;
    RECT 0 44.870 0.070 45.640 ;
    RECT 0 45.710 0.070 46.480 ;
    RECT 0 46.550 0.070 47.320 ;
    RECT 0 47.390 0.070 48.160 ;
    RECT 0 48.230 0.070 49.000 ;
    RECT 0 49.070 0.070 49.840 ;
    RECT 0 49.910 0.070 50.680 ;
    RECT 0 50.750 0.070 51.520 ;
    RECT 0 51.590 0.070 52.360 ;
    RECT 0 52.430 0.070 53.200 ;
    RECT 0 53.270 0.070 54.040 ;
    RECT 0 54.110 0.070 54.880 ;
    RECT 0 54.950 0.070 55.720 ;
    RECT 0 55.790 0.070 56.560 ;
    RECT 0 56.630 0.070 57.400 ;
    RECT 0 57.470 0.070 59.920 ;
    RECT 0 59.990 0.070 60.760 ;
    RECT 0 60.830 0.070 61.600 ;
    RECT 0 61.670 0.070 62.440 ;
    RECT 0 62.510 0.070 63.280 ;
    RECT 0 63.350 0.070 64.120 ;
    RECT 0 64.190 0.070 64.960 ;
    RECT 0 65.030 0.070 65.800 ;
    RECT 0 65.870 0.070 66.640 ;
    RECT 0 66.710 0.070 67.480 ;
    RECT 0 67.550 0.070 68.320 ;
    RECT 0 68.390 0.070 69.160 ;
    RECT 0 69.230 0.070 70.000 ;
    RECT 0 70.070 0.070 70.840 ;
    RECT 0 70.910 0.070 71.680 ;
    RECT 0 71.750 0.070 72.520 ;
    RECT 0 72.590 0.070 73.360 ;
    RECT 0 73.430 0.070 74.200 ;
    RECT 0 74.270 0.070 75.040 ;
    RECT 0 75.110 0.070 75.880 ;
    RECT 0 75.950 0.070 76.720 ;
    RECT 0 76.790 0.070 77.560 ;
    RECT 0 77.630 0.070 78.400 ;
    RECT 0 78.470 0.070 79.240 ;
    RECT 0 79.310 0.070 80.080 ;
    RECT 0 80.150 0.070 80.920 ;
    RECT 0 80.990 0.070 81.760 ;
    RECT 0 81.830 0.070 82.600 ;
    RECT 0 82.670 0.070 83.440 ;
    RECT 0 83.510 0.070 84.280 ;
    RECT 0 84.350 0.070 85.120 ;
    RECT 0 85.190 0.070 85.960 ;
    RECT 0 86.030 0.070 88.480 ;
    RECT 0 88.550 0.070 89.320 ;
    RECT 0 89.390 0.070 90.160 ;
    RECT 0 90.230 0.070 91.000 ;
    RECT 0 91.070 0.070 91.840 ;
    RECT 0 91.910 0.070 92.680 ;
    RECT 0 92.750 0.070 93.520 ;
    RECT 0 93.590 0.070 94.360 ;
    RECT 0 94.430 0.070 95.200 ;
    RECT 0 95.270 0.070 96.040 ;
    RECT 0 96.110 0.070 98.560 ;
    RECT 0 98.630 0.070 99.400 ;
    RECT 0 99.470 0.070 100.240 ;
    RECT 0 100.310 0.070 107.800 ;
    LAYER M17 ;
    RECT 0 0 152.190 2.800 ;
    RECT 0 105.000 152.190 107.800 ;
    RECT 0.000 2.800 2.660 105.000 ;
    RECT 2.940 2.800 4.900 105.000 ;
    RECT 5.180 2.800 7.140 105.000 ;
    RECT 7.420 2.800 9.380 105.000 ;
    RECT 9.660 2.800 11.620 105.000 ;
    RECT 11.900 2.800 13.860 105.000 ;
    RECT 14.140 2.800 16.100 105.000 ;
    RECT 16.380 2.800 18.340 105.000 ;
    RECT 18.620 2.800 20.580 105.000 ;
    RECT 20.860 2.800 22.820 105.000 ;
    RECT 23.100 2.800 25.060 105.000 ;
    RECT 25.340 2.800 27.300 105.000 ;
    RECT 27.580 2.800 29.540 105.000 ;
    RECT 29.820 2.800 31.780 105.000 ;
    RECT 32.060 2.800 34.020 105.000 ;
    RECT 34.300 2.800 36.260 105.000 ;
    RECT 36.540 2.800 38.500 105.000 ;
    RECT 38.780 2.800 40.740 105.000 ;
    RECT 41.020 2.800 42.980 105.000 ;
    RECT 43.260 2.800 45.220 105.000 ;
    RECT 45.500 2.800 47.460 105.000 ;
    RECT 47.740 2.800 49.700 105.000 ;
    RECT 49.980 2.800 51.940 105.000 ;
    RECT 52.220 2.800 54.180 105.000 ;
    RECT 54.460 2.800 56.420 105.000 ;
    RECT 56.700 2.800 58.660 105.000 ;
    RECT 58.940 2.800 60.900 105.000 ;
    RECT 61.180 2.800 63.140 105.000 ;
    RECT 63.420 2.800 65.380 105.000 ;
    RECT 65.660 2.800 67.620 105.000 ;
    RECT 67.900 2.800 69.860 105.000 ;
    RECT 70.140 2.800 72.100 105.000 ;
    RECT 72.380 2.800 74.340 105.000 ;
    RECT 74.620 2.800 76.580 105.000 ;
    RECT 76.860 2.800 78.820 105.000 ;
    RECT 79.100 2.800 81.060 105.000 ;
    RECT 81.340 2.800 83.300 105.000 ;
    RECT 83.580 2.800 85.540 105.000 ;
    RECT 85.820 2.800 87.780 105.000 ;
    RECT 88.060 2.800 90.020 105.000 ;
    RECT 90.300 2.800 92.260 105.000 ;
    RECT 92.540 2.800 94.500 105.000 ;
    RECT 94.780 2.800 96.740 105.000 ;
    RECT 97.020 2.800 98.980 105.000 ;
    RECT 99.260 2.800 101.220 105.000 ;
    RECT 101.500 2.800 103.460 105.000 ;
    RECT 103.740 2.800 105.700 105.000 ;
    RECT 105.980 2.800 107.940 105.000 ;
    RECT 108.220 2.800 110.180 105.000 ;
    RECT 110.460 2.800 112.420 105.000 ;
    RECT 112.700 2.800 114.660 105.000 ;
    RECT 114.940 2.800 116.900 105.000 ;
    RECT 117.180 2.800 119.140 105.000 ;
    RECT 119.420 2.800 121.380 105.000 ;
    RECT 121.660 2.800 123.620 105.000 ;
    RECT 123.900 2.800 125.860 105.000 ;
    RECT 126.140 2.800 128.100 105.000 ;
    RECT 128.380 2.800 130.340 105.000 ;
    RECT 130.620 2.800 132.580 105.000 ;
    RECT 132.860 2.800 134.820 105.000 ;
    RECT 135.100 2.800 137.060 105.000 ;
    RECT 137.340 2.800 139.300 105.000 ;
    RECT 139.580 2.800 141.540 105.000 ;
    RECT 141.820 2.800 143.780 105.000 ;
    RECT 144.060 2.800 146.020 105.000 ;
    RECT 146.300 2.800 148.260 105.000 ;
    RECT 148.540 2.800 152.190 105.000 ;
  END
END fakeram45_1024x32_upper

END LIBRARY
